#---------------------------------------------------------------------------#
# Text definition Poscalib.sv
# (c)Copyright ABB - 2004-09-28 15:32:09
#---------------------------------------------------------------------------#
#
Poscalib::
#
#
0: #tdrvIntrchCal
IRBP Stationsv�xel kalibrering
#
1: #tdrvStnCal
IRBP Station kalibrering
#
2: #tdrvIntCalStart
Starta kalibrering av stationsv�xel
#
3: #tdrvStnCalStart
Starta kalibrering av station
#
4: #tdrvCancelTxt
- Tryck Avbryt f�r att avsluta
#
5: #tdrvOKTxt
- Tryck OK f�r att forts�tta
#
6: #tdrvFkCancel
Avbryt
#
7: #tdrvFkOK
OK
#
8: #tdrvCalibFin
Kalibrering f�rdig.
#
9: #tdrvWrongOpMode
Fel k�rs�tt.
#
10: #tdrvOpModeMan
Tryck OK, �ndra till MANUELL
#
11: #tdrvOpModeManFs
Tryck OK, �ndra till MANUELL 100%
#
12: #tdrvOpModeAuto
Tryck OK, �ndra till AUTO
#
13: #tdrvOpModeRest
och starta om.
#
14: #tdrvRobMov1
F�rflytta roboten till en position
#
15: #tdrvRobMov2
d�r den kan st� medan kalib. p�g�r.
#
16: #tdrvRobMov3
Starta sedan om programmet.
#
17: #tdrvIntchMov1
Stationsv�xeln kan nu r�ra p� sig.
#
18: #tdrvIntchMov2
Se till att h�lla s�kerhetsavst�nd.
#
19: #tdrvIntchMov3
""
#
20: #tdrvIntchPos1
Stationsv�xeln �r inte i l�ge. Tryck
#
21: #tdrvIntchPos2
OK och jogga sedan stationsv�xeln
#
22: #tdrvIntchPos3
i position.
#
23: #tdrvCalDone1
Kalibrerar
#
24: #tdrvCalDone2
% f�rdigt...
#
25: #tdrvCalOkPr
1. Tryck OK.
#
26: #tdrvCalFine1
2. Finkalibrera
#
27: #tdrvCalFine2
axel
#
28: #tdrvCalRest
3. Starta om programmet.
#
29: #tdrvTorque
Moment:
#
30: #tdrvAngle
Vinkel:
#
31: #tdrvNM
(Nm)
#
32: #tdrvDeg
(deg)
#
33: #tdrvItchChk
IRBP stationsv�xel kontroll
#
34: #tdrvChkPos1
kontrollerar (sida 1)...
#
35: #tdrvChkPos2
kontrollerar (sida 2)...
#
36: #tdrvChkPos3
kontrollerar (sida 3)...
#
37: #tdrvChkPos4
kontrollerar (sida 4)...
#
38: #tdrvDataWrite
Data har skrivits fill fil.
#
39: #tdrvTPU
Ska data presenteras p� TPU?
#
40: #tdrvYES
Ja
#
41: #tdrvNO
Nej
#
42: #tdrvStnLA1
Sida 1. Vinkel 1=
#
43: #tdrvStnRA1
Sida 1. Vinkel 2=
#
44: #tdrvStnBA1
Sida 1. Brytvinkel=
#
45: #tdrvStnLA2
Sida 2. Vinkel 1=
#
46: #tdrvStnRA2
Sida 2. Vinkel 2=
#
47: #tdrvStnBA
Sida 2. Brytvinkel=
#
48: #tdrvStnLA3
Sida 3. Vinkel 1=
#
49: #tdrvStnRA3
Sida 3. Vinkel 2=
#
50: #tdrvStnBA3
Sida 3. Brytvinkel=
#
51: #tdrvStnLA4
Sida 4. Vinkel 1=
#
52: #tdrvStnRA4
Sida 4. Vinkel 2=
#
53: #tdrvStnBA4
Sida 4. Brytvinkel=
#
54: #tdrvTorqueErr1
F�r stort moment. Ta av last och
#
55: #tdrvTorqueErr2
k�r kalibrering igen.
#
56: #tdrvTorqueErr3
""
#
# END OF FILE
#
